/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Jan  3 07:38:57 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2088510296 */

module datapath(p_0, p_1);
   input [2:0]p_0;
   output [6:0]p_1;

   INV_X1 i_0 (.A(p_0[0]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[1]), .ZN(n_1));
   NAND2_X1 i_2 (.A1(n_0), .A2(n_1), .ZN(n_2));
   NAND2_X1 i_3 (.A1(p_0[0]), .A2(n_1), .ZN(n_3));
   NAND2_X1 i_4 (.A1(n_0), .A2(p_0[1]), .ZN(n_4));
   NAND2_X1 i_5 (.A1(p_0[0]), .A2(p_0[1]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NOR2_X1 i_7 (.A1(n_3), .A2(p_0[2]), .ZN(p_1[1]));
   NOR2_X1 i_8 (.A1(n_4), .A2(p_0[2]), .ZN(p_1[2]));
   NOR2_X1 i_9 (.A1(n_5), .A2(p_0[2]), .ZN(p_1[3]));
   NOR2_X1 i_10 (.A1(n_2), .A2(n_6), .ZN(p_1[4]));
   NOR2_X1 i_11 (.A1(n_3), .A2(n_6), .ZN(p_1[5]));
   NOR2_X1 i_12 (.A1(n_4), .A2(n_6), .ZN(p_1[6]));
endmodule

module FSMHomeAutomation(clk, rst, sensors, temp, output_signals, display);
   input clk;
   input rst;
   input [3:0]sensors;
   input [5:0]temp;
   output [5:0]output_signals;
   output [2:0]display;

   wire n_0_0;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_2_18;
   wire n_0_2_19;
   wire n_0_2_20;
   wire n_0_2_21;
   wire n_0_2_22;
   wire n_0_2_23;
   wire n_0_2_24;
   wire n_0_2_25;
   wire n_0_2_26;
   wire n_0_2_27;
   wire n_0_2_28;
   wire n_0_2_29;
   wire n_0_2_30;
   wire n_0_2_31;
   wire n_0_2_32;
   wire n_0_2_33;
   wire n_0_2_34;
   wire n_0_2_35;
   wire n_0_2_36;
   wire n_0_1;
   wire n_0_2_37;
   wire n_0_2_38;
   wire n_0_2_39;
   wire n_0_2_40;
   wire n_0_2_41;
   wire n_0_2_42;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_2_47;
   wire n_0_2_48;
   wire n_0_2_49;
   wire n_0_2_50;
   wire n_0_2_51;
   wire n_0_2_52;
   wire n_0_2_53;
   wire n_0_2_54;
   wire n_0_2_55;
   wire n_0_2_56;
   wire n_0_2_57;
   wire n_0_2_58;
   wire n_0_2_59;
   wire n_0_2_60;
   wire n_0_2_61;
   wire n_0_2_62;
   wire n_0_2_63;
   wire n_0_2_64;
   wire n_0_2_65;
   wire n_0_2_66;
   wire n_0_2_67;
   wire n_0_2_68;
   wire n_0_2_69;
   wire n_0_2_70;
   wire n_0_2;
   wire n_0_2_71;
   wire n_0_2_72;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_2_75;
   wire n_0_2_76;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_2_79;
   wire n_0_2_80;
   wire n_0_2_81;
   wire n_0_2_82;
   wire n_0_2_83;
   wire n_0_2_84;
   wire n_0_2_85;
   wire n_0_2_86;
   wire n_0_2_89;
   wire n_0_2_90;
   wire n_0_2_91;
   wire n_0_2_92;
   wire n_0_2_93;
   wire n_0_2_94;
   wire n_0_2_95;
   wire n_0_2_96;
   wire n_0_2_97;
   wire n_0_2_98;
   wire n_0_2_99;
   wire n_0_2_100;
   wire n_0_2_101;
   wire n_0_2_102;
   wire n_0_2_103;
   wire n_0_2_104;
   wire n_0_2_105;
   wire n_0_3;
   wire n_0_2_87;
   wire n_0_2_88;
   wire n_0_3_0;
   wire n_0_3_1;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_4_0;
   wire n_0_13;
   wire n_0_4_1;
   wire n_0_4_2;
   wire n_0_4_3;
   wire n_0_4_4;
   wire n_0_4_5;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;

   DFF_X1 \currentstate_reg[2]  (.D(n_0_12), .CK(clk), .Q(display[2]), .QN());
   DFF_X1 \currentstate_reg[1]  (.D(n_0_11), .CK(clk), .Q(display[1]), .QN());
   DFF_X1 \currentstate_reg[0]  (.D(n_0_10), .CK(clk), .Q(display[0]), .QN());
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(n_0_0));
   NAND2_X1 i_0_0_1 (.A1(n_0_0_5), .A2(n_0_0_1), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_2), .ZN(n_0_0_1));
   NAND2_X1 i_0_0_3 (.A1(n_0_0_4), .A2(n_0_0_3), .ZN(n_0_0_2));
   INV_X1 i_0_0_4 (.A(temp[4]), .ZN(n_0_0_3));
   INV_X1 i_0_0_5 (.A(temp[5]), .ZN(n_0_0_4));
   OAI21_X1 i_0_0_6 (.A(temp[3]), .B1(temp[2]), .B2(temp[1]), .ZN(n_0_0_5));
   NAND2_X1 i_0_2_0 (.A1(n_0_13), .A2(n_0_2_52), .ZN(n_0_2_0));
   NAND3_X1 i_0_2_1 (.A1(n_0_2_61), .A2(n_0_2_79), .A3(n_0_2_54), .ZN(n_0_2_1));
   NAND2_X1 i_0_2_2 (.A1(n_0_2_71), .A2(display[1]), .ZN(n_0_2_2));
   NOR2_X1 i_0_2_3 (.A1(n_0_2_55), .A2(n_0_2_2), .ZN(n_0_2_3));
   NAND2_X1 i_0_2_4 (.A1(n_0_2_61), .A2(n_0_2_3), .ZN(n_0_2_4));
   INV_X1 i_0_2_5 (.A(n_0_2_51), .ZN(n_0_2_5));
   NAND2_X1 i_0_2_6 (.A1(n_0_2_5), .A2(n_0_2_37), .ZN(n_0_2_6));
   NAND3_X1 i_0_2_7 (.A1(n_0_2_1), .A2(n_0_2_4), .A3(n_0_2_6), .ZN(n_0_2_7));
   NAND3_X1 i_0_2_8 (.A1(n_0_2_0), .A2(n_0_0), .A3(n_0_2_7), .ZN(n_0_2_8));
   NOR2_X1 i_0_2_9 (.A1(n_0_2_2), .A2(display[0]), .ZN(n_0_2_9));
   OAI22_X1 i_0_2_10 (.A1(n_0_2_76), .A2(display[0]), .B1(display[2]), .B2(
      display[1]), .ZN(n_0_2_10));
   NOR2_X1 i_0_2_11 (.A1(n_0_2_9), .A2(n_0_2_10), .ZN(n_0_2_11));
   INV_X1 i_0_2_12 (.A(n_0_2_11), .ZN(n_0_2_12));
   NAND3_X1 i_0_2_13 (.A1(n_0_2_79), .A2(sensors[2]), .A3(n_0_2_12), .ZN(
      n_0_2_13));
   INV_X1 i_0_2_14 (.A(n_0_2_2), .ZN(n_0_2_14));
   NAND2_X1 i_0_2_15 (.A1(n_0_2_14), .A2(n_0_2_37), .ZN(n_0_2_15));
   NOR2_X1 i_0_2_16 (.A1(n_0_2_11), .A2(n_0_2_15), .ZN(n_0_2_16));
   NAND2_X1 i_0_2_17 (.A1(sensors[2]), .A2(n_0_2_16), .ZN(n_0_2_17));
   XNOR2_X1 i_0_2_18 (.A(display[2]), .B(display[1]), .ZN(n_0_2_18));
   NAND2_X1 i_0_2_19 (.A1(n_0_2_18), .A2(n_0_2_37), .ZN(n_0_2_19));
   INV_X1 i_0_2_20 (.A(n_0_2_19), .ZN(n_0_2_20));
   NAND2_X1 i_0_2_21 (.A1(sensors[0]), .A2(n_0_2_20), .ZN(n_0_2_21));
   NAND3_X1 i_0_2_22 (.A1(n_0_2_13), .A2(n_0_2_17), .A3(n_0_2_21), .ZN(n_0_2_22));
   INV_X1 i_0_2_23 (.A(n_0_13), .ZN(n_0_2_23));
   NAND2_X1 i_0_2_24 (.A1(n_0_2_83), .A2(n_0_2_2), .ZN(n_0_2_24));
   NAND3_X1 i_0_2_25 (.A1(n_0_2_61), .A2(n_0_2_79), .A3(n_0_2_24), .ZN(n_0_2_25));
   NAND2_X1 i_0_2_26 (.A1(n_0_2_24), .A2(n_0_2_77), .ZN(n_0_2_26));
   INV_X1 i_0_2_27 (.A(n_0_2_26), .ZN(n_0_2_27));
   NAND2_X1 i_0_2_28 (.A1(n_0_2_61), .A2(n_0_2_27), .ZN(n_0_2_28));
   NAND2_X1 i_0_2_29 (.A1(n_0_2_24), .A2(n_0_2_37), .ZN(n_0_2_29));
   INV_X1 i_0_2_30 (.A(n_0_2_29), .ZN(n_0_2_30));
   NAND2_X1 i_0_2_31 (.A1(n_0_2_61), .A2(n_0_2_30), .ZN(n_0_2_31));
   NAND4_X1 i_0_2_32 (.A1(n_0_2_25), .A2(n_0_2_28), .A3(n_0_2_31), .A4(n_0_2_51), 
      .ZN(n_0_2_32));
   OAI21_X1 i_0_2_33 (.A(n_0_2_80), .B1(n_0_2_75), .B2(sensors[1]), .ZN(n_0_2_33));
   NAND2_X1 i_0_2_34 (.A1(n_0_2_32), .A2(n_0_2_33), .ZN(n_0_2_34));
   INV_X1 i_0_2_35 (.A(n_0_2_34), .ZN(n_0_2_35));
   AOI21_X1 i_0_2_36 (.A(n_0_2_22), .B1(n_0_2_23), .B2(n_0_2_35), .ZN(n_0_2_36));
   NAND2_X1 i_0_2_37 (.A1(n_0_2_8), .A2(n_0_2_36), .ZN(n_0_1));
   INV_X1 i_0_2_38 (.A(display[0]), .ZN(n_0_2_37));
   NAND3_X1 i_0_2_39 (.A1(n_0_2_37), .A2(n_0_2_71), .A3(display[1]), .ZN(
      n_0_2_38));
   NAND2_X1 i_0_2_40 (.A1(sensors[1]), .A2(n_0_2_38), .ZN(n_0_2_39));
   NAND2_X1 i_0_2_41 (.A1(n_0_2_39), .A2(n_0_2_75), .ZN(n_0_2_40));
   XNOR2_X1 i_0_2_42 (.A(display[0]), .B(display[1]), .ZN(n_0_2_41));
   INV_X1 i_0_2_43 (.A(n_0_2_41), .ZN(n_0_2_42));
   NAND2_X1 i_0_2_44 (.A1(n_0_2_42), .A2(n_0_2_71), .ZN(n_0_2_43));
   NAND2_X1 i_0_2_45 (.A1(sensors[0]), .A2(n_0_2_43), .ZN(n_0_2_44));
   NAND2_X1 i_0_2_46 (.A1(n_0_2_71), .A2(n_0_2_76), .ZN(n_0_2_45));
   NAND2_X1 i_0_2_47 (.A1(n_0_2_41), .A2(n_0_2_45), .ZN(n_0_2_46));
   INV_X1 i_0_2_48 (.A(n_0_2_46), .ZN(n_0_2_47));
   NAND2_X1 i_0_2_49 (.A1(n_0_2_43), .A2(n_0_2_47), .ZN(n_0_2_48));
   NAND3_X1 i_0_2_50 (.A1(n_0_2_40), .A2(n_0_2_44), .A3(n_0_2_48), .ZN(n_0_2_49));
   INV_X1 i_0_2_51 (.A(n_0_2_49), .ZN(n_0_2_50));
   NAND2_X1 i_0_2_52 (.A1(n_0_2_76), .A2(display[2]), .ZN(n_0_2_51));
   NOR2_X1 i_0_2_53 (.A1(n_0_2_51), .A2(n_0_2_37), .ZN(n_0_2_52));
   AOI21_X1 i_0_2_54 (.A(n_0_2_50), .B1(n_0_13), .B2(n_0_2_52), .ZN(n_0_2_53));
   NAND3_X1 i_0_2_55 (.A1(display[0]), .A2(display[2]), .A3(display[1]), 
      .ZN(n_0_2_54));
   INV_X1 i_0_2_56 (.A(n_0_2_54), .ZN(n_0_2_55));
   NOR2_X1 i_0_2_57 (.A1(sensors[0]), .A2(n_0_2_55), .ZN(n_0_2_56));
   NAND2_X1 i_0_2_58 (.A1(n_0_2_75), .A2(n_0_2_79), .ZN(n_0_2_57));
   NAND2_X1 i_0_2_59 (.A1(sensors[3]), .A2(display[1]), .ZN(n_0_2_58));
   NAND3_X1 i_0_2_60 (.A1(n_0_2_56), .A2(n_0_2_57), .A3(n_0_2_58), .ZN(n_0_2_59));
   INV_X1 i_0_2_61 (.A(n_0_2_59), .ZN(n_0_2_60));
   INV_X1 i_0_2_62 (.A(sensors[3]), .ZN(n_0_2_61));
   OAI21_X1 i_0_2_63 (.A(display[0]), .B1(n_0_2_98), .B2(display[2]), .ZN(
      n_0_2_62));
   NAND3_X1 i_0_2_64 (.A1(n_0_2_61), .A2(n_0_2_80), .A3(n_0_2_62), .ZN(n_0_2_63));
   INV_X1 i_0_2_65 (.A(n_0_2_62), .ZN(n_0_2_64));
   INV_X1 i_0_2_66 (.A(n_0_2_98), .ZN(n_0_2_65));
   NAND2_X1 i_0_2_67 (.A1(n_0_2_65), .A2(n_0_2_71), .ZN(n_0_2_66));
   NOR2_X1 i_0_2_68 (.A1(n_0_2_64), .A2(n_0_2_66), .ZN(n_0_2_67));
   NAND2_X1 i_0_2_69 (.A1(n_0_2_61), .A2(n_0_2_67), .ZN(n_0_2_68));
   NAND3_X1 i_0_2_70 (.A1(n_0_2_63), .A2(n_0_2_68), .A3(n_0_2_51), .ZN(n_0_2_69));
   AOI21_X1 i_0_2_71 (.A(n_0_2_60), .B1(n_0_13), .B2(n_0_2_69), .ZN(n_0_2_70));
   OAI21_X1 i_0_2_72 (.A(n_0_2_53), .B1(n_0_2_70), .B2(n_0_0), .ZN(n_0_2));
   INV_X1 i_0_2_73 (.A(display[2]), .ZN(n_0_2_71));
   NAND2_X1 i_0_2_74 (.A1(n_0_2_71), .A2(display[0]), .ZN(n_0_2_72));
   INV_X1 i_0_2_75 (.A(n_0_2_72), .ZN(n_0_2_73));
   MUX2_X1 i_0_2_76 (.A(display[2]), .B(n_0_2_73), .S(display[1]), .Z(n_0_2_74));
   INV_X1 i_0_2_77 (.A(sensors[2]), .ZN(n_0_2_75));
   INV_X1 i_0_2_78 (.A(display[1]), .ZN(n_0_2_76));
   NOR2_X1 i_0_2_79 (.A1(n_0_2_76), .A2(display[2]), .ZN(n_0_2_77));
   AOI21_X1 i_0_2_80 (.A(n_0_2_74), .B1(n_0_2_75), .B2(n_0_2_77), .ZN(n_0_2_78));
   INV_X1 i_0_2_81 (.A(sensors[1]), .ZN(n_0_2_79));
   INV_X1 i_0_2_82 (.A(sensors[0]), .ZN(n_0_2_80));
   NAND2_X1 i_0_2_83 (.A1(display[0]), .A2(display[1]), .ZN(n_0_2_81));
   NAND4_X1 i_0_2_84 (.A1(n_0_2_79), .A2(n_0_2_80), .A3(n_0_2_75), .A4(n_0_2_81), 
      .ZN(n_0_2_82));
   INV_X1 i_0_2_85 (.A(n_0_2_81), .ZN(n_0_2_83));
   NAND2_X1 i_0_2_86 (.A1(n_0_2_76), .A2(display[0]), .ZN(n_0_2_84));
   NOR2_X1 i_0_2_87 (.A1(n_0_2_83), .A2(n_0_2_84), .ZN(n_0_2_85));
   NAND3_X1 i_0_2_88 (.A1(n_0_2_79), .A2(n_0_2_75), .A3(n_0_2_85), .ZN(n_0_2_86));
   NAND3_X1 i_0_2_91 (.A1(n_0_2_76), .A2(display[0]), .A3(display[2]), .ZN(
      n_0_2_89));
   INV_X1 i_0_2_92 (.A(n_0_2_89), .ZN(n_0_2_90));
   NAND2_X1 i_0_2_93 (.A1(sensors[2]), .A2(n_0_2_90), .ZN(n_0_2_91));
   NAND2_X1 i_0_2_94 (.A1(sensors[0]), .A2(n_0_2_90), .ZN(n_0_2_92));
   NAND2_X1 i_0_2_95 (.A1(sensors[1]), .A2(n_0_2_90), .ZN(n_0_2_93));
   NAND3_X1 i_0_2_96 (.A1(n_0_2_91), .A2(n_0_2_92), .A3(n_0_2_93), .ZN(n_0_2_94));
   INV_X1 i_0_2_97 (.A(n_0_2_94), .ZN(n_0_2_95));
   NAND2_X1 i_0_2_98 (.A1(n_0_0), .A2(n_0_2_95), .ZN(n_0_2_96));
   NAND3_X1 i_0_2_99 (.A1(n_0_2_92), .A2(n_0_2_93), .A3(sensors[3]), .ZN(
      n_0_2_97));
   NOR2_X1 i_0_2_100 (.A1(display[0]), .A2(display[1]), .ZN(n_0_2_98));
   NAND2_X1 i_0_2_101 (.A1(sensors[2]), .A2(n_0_2_98), .ZN(n_0_2_99));
   NAND2_X1 i_0_2_102 (.A1(sensors[0]), .A2(n_0_2_98), .ZN(n_0_2_100));
   NAND2_X1 i_0_2_103 (.A1(n_0_2_99), .A2(n_0_2_100), .ZN(n_0_2_101));
   NAND2_X1 i_0_2_104 (.A1(sensors[1]), .A2(n_0_2_98), .ZN(n_0_2_102));
   NAND2_X1 i_0_2_105 (.A1(n_0_2_102), .A2(n_0_2_91), .ZN(n_0_2_103));
   NOR3_X1 i_0_2_106 (.A1(n_0_2_97), .A2(n_0_2_101), .A3(n_0_2_103), .ZN(
      n_0_2_104));
   NOR2_X1 i_0_2_107 (.A1(n_0_13), .A2(n_0_2_104), .ZN(n_0_2_105));
   AOI21_X1 i_0_2_108 (.A(n_0_2_88), .B1(n_0_2_96), .B2(n_0_2_105), .ZN(n_0_3));
   NAND3_X1 i_0_2_89 (.A1(n_0_2_82), .A2(n_0_2_86), .A3(n_0_2_78), .ZN(n_0_2_87));
   INV_X1 i_0_2_90 (.A(n_0_2_87), .ZN(n_0_2_88));
   INV_X1 i_0_3_0 (.A(rst), .ZN(n_0_3_0));
   NAND3_X1 i_0_3_1 (.A1(n_0_3), .A2(n_0_2), .A3(n_0_1), .ZN(n_0_3_1));
   AND3_X1 i_0_3_2 (.A1(n_0_14), .A2(n_0_3_0), .A3(n_0_3_1), .ZN(n_0_4));
   AND3_X1 i_0_3_3 (.A1(n_0_15), .A2(n_0_3_1), .A3(n_0_3_0), .ZN(n_0_5));
   AND3_X1 i_0_3_4 (.A1(n_0_3_1), .A2(n_0_16), .A3(n_0_3_0), .ZN(n_0_6));
   AND3_X1 i_0_3_5 (.A1(n_0_17), .A2(n_0_3_0), .A3(n_0_3_1), .ZN(n_0_7));
   AND3_X1 i_0_3_6 (.A1(n_0_18), .A2(n_0_3_0), .A3(n_0_3_1), .ZN(n_0_8));
   AND3_X1 i_0_3_7 (.A1(n_0_19), .A2(n_0_3_0), .A3(n_0_3_1), .ZN(n_0_9));
   AND2_X1 i_0_4_0 (.A1(n_0_4_0), .A2(n_0_1), .ZN(n_0_10));
   AND2_X1 i_0_4_1 (.A1(n_0_4_0), .A2(n_0_2), .ZN(n_0_11));
   AND2_X1 i_0_4_2 (.A1(n_0_4_0), .A2(n_0_3), .ZN(n_0_12));
   INV_X1 i_0_4_3 (.A(rst), .ZN(n_0_4_0));
   NAND2_X1 i_0_4_4 (.A1(n_0_4_1), .A2(n_0_4_5), .ZN(n_0_13));
   NAND2_X1 i_0_4_5 (.A1(n_0_4_2), .A2(temp[4]), .ZN(n_0_4_1));
   NAND2_X1 i_0_4_6 (.A1(n_0_4_3), .A2(n_0_4_4), .ZN(n_0_4_2));
   NAND2_X1 i_0_4_7 (.A1(temp[2]), .A2(temp[1]), .ZN(n_0_4_3));
   INV_X1 i_0_4_8 (.A(temp[3]), .ZN(n_0_4_4));
   INV_X1 i_0_4_9 (.A(temp[5]), .ZN(n_0_4_5));
   datapath i_0_1 (.p_0({n_0_3, n_0_2, n_0_1}), .p_1({n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, uc_0}));
   DFF_X2 \temp_output_signals_reg[2]  (.D(n_0_6), .CK(clk), .Q(
      output_signals[2]), .QN());
   DFF_X1 \temp_output_signals_reg[1]  (.D(n_0_5), .CK(clk), .Q(
      output_signals[1]), .QN());
   DFF_X1 \temp_output_signals_reg[5]  (.D(n_0_9), .CK(clk), .Q(
      output_signals[5]), .QN());
   DFF_X1 \temp_output_signals_reg[3]  (.D(n_0_7), .CK(clk), .Q(
      output_signals[3]), .QN());
   DFF_X1 \temp_output_signals_reg[4]  (.D(n_0_8), .CK(clk), .Q(
      output_signals[4]), .QN());
   DFF_X1 \temp_output_signals_reg[0]  (.D(n_0_4), .CK(clk), .Q(
      output_signals[0]), .QN());
endmodule
